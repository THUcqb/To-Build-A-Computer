----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    20:57:08 11/09/2017
-- Design Name:
-- Module Name:    MemoryAndSerialPort - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MemoryAndSerialPort is
end MemoryAndSerialPort;

architecture Behavioral of MemoryAndSerialPort is

begin


end Behavioral;

